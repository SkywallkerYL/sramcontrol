`ifndef macro__SV
`define macro__SV

`define SimulationTime 1400000

`define readTime 70000

`define itemnum 10

`endif