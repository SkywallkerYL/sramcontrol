`ifndef MY_MONITOR__SV
`define MY_MONITOR__SV
class my_monitor extends uvm_monitor;

   virtual fiforead_if vif;

   uvm_analysis_port #(my_transaction)  ap;
   
   `uvm_component_utils(my_monitor)
   function new(string name = "my_monitor", uvm_component parent = null);
      super.new(name, parent);
   endfunction

   virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      if(!uvm_config_db#(virtual fiforead_if)::get(this, "", "vif", vif))
         `uvm_fatal("my_monitor", "virtual interface must be set for vif!!!")
      ap = new("ap", this);
   endfunction

   extern task main_phase(uvm_phase phase);
   extern task collect_one_pkt(my_transaction tr);
endclass

task my_monitor::main_phase(uvm_phase phase);
   my_transaction tr;
   while(1) begin
      tr = new("tr");
      collect_one_pkt(tr);
      //tr.print();
      ap.write(tr);
   end
endtask

task my_monitor::collect_one_pkt(my_transaction tr);
   byte unsigned data_q[$];
   byte unsigned data_array[];
   logic [15:0] data;
   logic readen = 0;
   logic empty = 0;
   int data_size;
   
   while(1) begin
      @(posedge vif.rclk);
      if(!vif.empty) break;
   end
   
   `uvm_info("my_monitor", "begin to collect one pkt", UVM_LOW);
   vif.readen <= 1'b1;
   @(posedge vif.rclk);
  
   //while(!vif.empty) begin
      @(posedge vif.rclk);
      data_q.push_back(vif.data);
      $display("monitor data: %d",vif.data);
      vif.readen <= 1'b0;
      @(posedge vif.rclk); 
      
      data_q.push_back(vif.data);
      $display("monitor data: %d",vif.data);
      //@(posedge vif.rclk);
   //end
   data_size  = data_q.size();   
   data_array = new[data_size];
   for ( int i = 0; i < data_size; i++ ) begin
      data_array[i] = data_q[i];
      
      //tr.print(data);
   end
   
   //这里使用unpack_bytes函数将data_q中的byte流转换成tr中的各个字段。unpack_bytes函数的输入参数必须是一个动态数组，所
//以需要先把收集到的、放在data_q中的数据复制到一个动态数组中。由于tr中的pload是一个动态数组，所以需要在调用
//unpack_bytes之前指定其大小，这样unpack_bytes函数才能正常工作。
   //tr.pload = new[data_size - 18]; //da sa, e_type, crc
   data_size = tr.unpack_bytes(data_array) / 8; 
   //tr.print();
   `uvm_info("my_monitor", "end collect one pkt", UVM_LOW);
endtask


`endif
