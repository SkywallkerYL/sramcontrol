`ifndef macro__SV
`define macro__SV

`define SimulationTime 100000

`define readTime 50000

`define itemnum 10


`endif